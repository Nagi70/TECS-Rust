import("struct.cdl");
import("time_delay_kalman_filter.cdl");
import("state_transition.cdl");
import("measurement.cdl");
import("mahalanobis.cdl");
import("covariance.cdl");
import("utils_geometry.cdl");

signature sEkfModule {
    void init( void );
    void accumulateDelayTime( [in] double64_t dt );
    int32_t findClosestDelayTimeIndex( [in] double64_t target_value); // measurementUpdateTwist に埋め込む方がいいかも
    void predictWithDelay([in] double64_t dt );
    PLType("Result<(), EkfModuleError>") measurementUpdateTwist( [in] struct TwistWithCovariance twist, [in] PLTYpe("awkernel_lib::time::Time") ccurent_time );　// エラーenumはユーザ定義
    void getCurrentTwist( [in] PLTYpe("awkernel_lib::time::Time") ccurent_time, [out] struct TwistWithCovarianceStamped* twist );
    void getCurrentTwistCovariance( [out] struct TwistWithCovariance twist );
    void getCurrentPoseCovariance( [out] struct PoseWithCovariance pose );
};

struct Simple1DFilter {
    double64_t x;
    double64_t var;
};

[generate( RustAWKPlugin , "")]
celltype tEkfModule {
    call sTimeDelayKalmanFilter     cKalman;
    call sStateTransition           cState;
    call sMeasurement               cMeasure;
    call sMahalanobis               cMaha;
    call sCovariance                cCov;
    call sUtilsGeometry             cUtils;

    entry sEkfModule eEkfModule;

    attr {
        int32_t extend_state_step = 50;
        bool_t enable_yaw_bias_estimation = true;

        double64_t z_filter_proc_dev = 5.0;
        double64_t roll_filter_proc_dev = 0.1;
        double64_t pitch_filter_proc_dev = 0.1;

        double64_t proc_stddev_yaw_c = 0.005;
        double64_t proc_stddev_vx_c = 10.0;
        double64_t proc_stddev_wz_c = 5.0;

        int32_t dim_x = 6;

        /* twistゲート・平滑化 */
        double64_t  twist_gate_dist = 46.1;
        uint32_t twist_smoothing_steps = 2;
        double64_t  twist_additional_delay = 0.0;

        // 初期位置情報 (下記のtfをあらかじめ加味してもいい)
        struct PoseWithCovariance initial_pose = {
            {
                PL_EXP("nalgebra::Vector3::new(1, 1, 1)"),
                PL_EXP("nalgebra::Quaternion::new(1, 2, 3, 4)")
            },
            PL_EXP("nalgebra::Matrix6::new(
                1, 1, 1, 1, 1, 1,
                1, 1, 1, 1, 1, 1,
                1, 1, 1, 1, 1, 1,
                1, 1, 1, 1, 1, 1,
                1, 1, 1, 1, 1, 1,
                1, 1, 1, 1, 1, 1 )"
            )
        };

        // mapへの変換tf (マップと初期位置が固定ならおそらくTFも固定)
        struct Transform tf = {
            PL_EXP("nalgebra::Vector3::new(1, 1, 1)"),
            PL_EXP("nalgebra::Quaternion::new(1, 2, 3, 4)")
        };
    };

    var {
        [size_is(extend_state_step)]
        double64_t *accumulated_delay_times = {};
        double ekf_dt;
        /* DRでは角速度の履歴だけ最小保持（必要に応じて） */
        PLType("nalgebra::Vector3<f64>") last_angular_velocity;
        struct Simple1DFilter z_filter = {0.0, 0.0};
        struct Simple1DFilter roll_filter = {0.0, 0.0};
        struct Simple1DFilter pitch_filter = {0.0, 0.0};
    };
};
