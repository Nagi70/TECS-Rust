/*
 *  TOPPERS/ASP Kernel
 *      Toyohashi Open Platform for Embedded Real-Time Systems/
 *      Advanced Standard Profile Kernel
 * 
 *  Copyright (C) 2015,2016 by Ushio Laboratory
 *              Graduate School of Engineering Science, Osaka Univ., JAPAN
 *  Copyright (C) 2015-2020 by Embedded and Real-Time Systems Laboratory
 *              Graduate School of Information Science, Nagoya Univ., JAPAN
 * 
 *  上記著作権者は，以下の(1)〜(4)の条件を満たす場合に限り，本ソフトウェ
 *  ア（本ソフトウェアを改変したものを含む．以下同じ）を使用・複製・改
 *  変・再配布（以下，利用と呼ぶ）することを無償で許諾する．
 *  (1) 本ソフトウェアをソースコードの形で利用する場合には，上記の著作
 *      権表示，この利用条件および下記の無保証規定が，そのままの形でソー
 *      スコード中に含まれていること．
 *  (2) 本ソフトウェアを，ライブラリ形式など，他のソフトウェア開発に使
 *      用できる形で再配布する場合には，再配布に伴うドキュメント（利用
 *      者マニュアルなど）に，上記の著作権表示，この利用条件および下記
 *      の無保証規定を掲載すること．
 *  (3) 本ソフトウェアを，機器に組み込むなど，他のソフトウェア開発に使
 *      用できない形で再配布する場合には，次のいずれかの条件を満たすこ
 *      と．
 *    (a) 再配布に伴うドキュメント（利用者マニュアルなど）に，上記の著
 *        作権表示，この利用条件および下記の無保証規定を掲載すること．
 *    (b) 再配布の形態を，別に定める方法によって，TOPPERSプロジェクトに
 *        報告すること．
 *  (4) 本ソフトウェアの利用により直接的または間接的に生じるいかなる損
 *      害からも，上記著作権者およびTOPPERSプロジェクトを免責すること．
 *      また，本ソフトウェアのユーザまたはエンドユーザからのいかなる理
 *      由に基づく請求からも，上記著作権者およびTOPPERSプロジェクトを
 *      免責すること．
 * 
 *  本ソフトウェアは，無保証で提供されているものである．上記著作権者お
 *  よびTOPPERSプロジェクトは，本ソフトウェアに関して，特定の使用目的
 *  に対する適合性も含めて，いかなる保証も行わない．また，本ソフトウェ
 *  アの利用により直接的または間接的に生じたいかなる損害に関しても，そ
 *  の責任を負わない．
 * 
 *  $Id: kernel.cdl 1437 2020-05-20 12:12:16Z ertl-hiro $
 */

/*
 *		TOPPERS/ASPカーネルオブジェクト コンポーネント記述ファイル
 */

/*
 *  カーネルオブジェクトのコンポーネント化のためのヘッダファイル
 */
import_C("tecs_kernel.h");

typedef	int_t	TaskRef;

/*
 *  タスク本体のシグニチャ
 */
signature sTaskBody {
	void	main(void);
};

/*
 *  タスク操作のシグニチャ（タスクコンテキスト用）
 */
signature sTask {
	ER		activate(void);
	ER_UINT	cancelActivate(void);
	ER		getTaskState([out] STAT *p_tskstat);
	ER		changePriority([in] PRI priority);
	ER		getPriority([out] PRI *p_priority);
	ER		refer([out] T_RTSK *pk_taskStatus);

	ER		wakeup(void);
	ER_UINT	cancelWakeup(void);
	ER		releaseWait(void);
	ER		suspend(void);
	ER		resume(void);

	ER		raiseTerminate(void);
	ER		terminate(void);
};

/*
 *  タスク操作のシグニチャ（非タスクコンテキスト用）
 */
[context("non-task")]
signature siTask {
	ER		activate(void);
	ER		wakeup(void);
	ER		releaseWait(void);
};

/*
 *  タイムイベント通知を受け取るためのシグネチャ
 */
[context("non-task")]
signature siNotificationHandler {
};

/*
 *  タスクのセルタイプ
 */
[active, generate( RustASP3Plugin, "lib, TASK")]
celltype tTaskRs {
	[inline] entry	sTask	eTask;
	[inline] entry	siTask	eiTask;
	call	sTaskBody	cTaskBody;

	[inline] entry	siNotificationHandler	eiActivateNotificationHandler;
	[inline] entry	siNotificationHandler	eiWakeUpNotificationHandler;

	attr {
		[omit]ID		id = C_EXP("TECS_RUST_TASK$id$");
		//TaskRef			task = C_EXP("TSKID_$id$_REF");
		TaskRef			task_ref = C_EXP("unsafe{TaskRef::from_raw_nonnull(NonZeroI32::new(TECS_RUST_TASK$id$).unwrap())}");
		[omit] ATR		attribute = C_EXP("TA_NULL");
		[omit] PRI		priority;
		[omit] size_t	stackSize;
	};

	factory {
		//write("tecsgen.cfg",
		//		"CRE_TSK(%s, { %s, 0, tTask_start, %s, %s, NULL });",
		//							id, attribute, priority, stackSize);
		//write("kernel_obj_ref.rs", 
		//		"static %s_REF:TaskRef = unsafe{TaskRef::from_raw_nonnull(NonZeroI32::new(%s).unwrap())};",
		//							id, id);

	};
	FACTORY {
		//write("tecsgen.cfg", "#include \"$ct$_tecsgen.h\"");
		//write("$ct$_factory.h", "#include \"kernel_cfg.h\"");
		//write("lib.rs", "mod kernel_cfg;");
		//write("lib.rs", "mod kernel_obj_ref;");
		//write("kernel_obj_ref.rs", "use crate::kernel_cfg::*;");
	};
};
