const int32_t DIM_X = 6;
const int32_t DIM_Y_TWIST = 2;
const int32_t DIM_X_EX = 300;