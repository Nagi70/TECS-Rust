import("struct_define.cdl");

signature sImuRaw {
};

signature sImuData {
};

signature sImu {
};