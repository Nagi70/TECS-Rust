//typedef uint32_t Cow;
//typedef uint32_t SchedulerType;
//typedef uint32_t Duration;

//*** リアクター共通シグニチャ ***//
signature sReactorbody {
    void main(void);
};

//*** 周期リアクターセルタイプ ***//
[active, generate( RustAWKPlugin, "DAG_PERIODIC_REACTOR")]
celltype tDagPeriodicReactor {
    call sReactorbody cDagPeriodicReactorbody;
    //entry sTask eTask;
    
    attr{
        [omit] RType("Cow") name = PL_EXP("task_id");
        [omit] RType("Cow") publishTopicNames = PL_EXP("Topic1, Topic2");
        [omit] RType("SchedulerType") schedType = PL_EXP("SchedulerType::PrioritizedFIFO(7)");
        [omit] RType("Duration") period = PL_EXP("Duration::from_secs(1)");
    };
};

//*** 通常リアクターセルタイプ ***//
[active, generate( RustAWKPlugin, "DAG_REACTOR")]
celltype tDagReactor {
    call sReactorbody cDagReactorbody;
    //entry sTask eTask;
    
    attr{
        [omit] RType("Cow") name = PL_EXP("task_id");
        [omit] RType("Cow") subscribeTopicNames = PL_EXP("Topic1, Topic2");
        [omit] RType("Cow") publishTopicNames = PL_EXP("Topic3, Topic4");
        [omit] RType("SchedulerType") schedType = PL_EXP("SchedulerType::PrioritizedFIFO(7)");
    };
};

//*** シンクリアクターセルタイプ ***//
[active, generate( RustAWKPlugin, "DAG_SINK_REACTOR")]
celltype tDagSinkReactor {
    call sReactorbody cDagSinkReactorbody;
    //entry sTask eTask;
    
    attr{
        [omit] RType("Cow") name = PL_EXP("task_id");
        [omit] RType("Cow") subscribeTopicNames = PL_EXP("Topic3, Topic4");
        [omit] RType("SchedulerType") schedType = PL_EXP("SchedulerType::PrioritizedFIFO(7)");
        [omit] RType("Duration") relative_deadline = PL_EXP("Duration::from_secs(1)");
    };
};

//*** 周期リアクターセルタイプ ***//
[active, generate( RustAWKPlugin, "PERIODIC_REACTOR")]
celltype tPeriodicReactor {
    call sReactorbody cPeriodicReactorbody;
    //entry sTask eTask;
    
    attr{
        [omit] RType("Cow") name = PL_EXP("task_id");
        [omit] RType("Cow") publishTopicNames = PL_EXP("Topic1, Topic2");
        [omit] RType("SchedulerType") schedType = PL_EXP("SchedulerType::PrioritizedFIFO(7)");
        [omit] RType("Duration") period = PL_EXP("Duration::from_secs(1)");
    };
};

//*** 通常リアクターセルタイプ ***//
[active, generate( RustAWKPlugin, "REACTOR")]
celltype tReactor {
    call sReactorbody cReactorbody;
    //entry sTask eTask;
    
    attr{
        [omit] RType("Cow") name = PL_EXP("task_id");
        [omit] RType("Cow") subscribeTopicNames = PL_EXP("Topic1, Topic2");
        [omit] RType("Cow") publishTopicNames = PL_EXP("Topic3, Topic4");
        [omit] RType("SchedulerType") schedType = PL_EXP("SchedulerType::PrioritizedFIFO(7)");
    };
};

//*** シンクリアクターセルタイプ ***//
[active, generate( RustAWKPlugin, "SINK_REACTOR")]
celltype tSinkReactor {
    call sReactorbody cSinkReactorbody;
    //entry sTask eTask;
    
    attr{
        [omit] RType("Cow") name = PL_EXP("task_id");
        [omit] RType("Cow") subscribeTopicNames = PL_EXP("Topic3, Topic4");
        [omit] RType("SchedulerType") schedType = PL_EXP("SchedulerType::PrioritizedFIFO(7)");
        [omit] RType("Duration") relative_deadline = PL_EXP("Duration::from_secs(1)");
    };
};