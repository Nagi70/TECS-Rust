signature sUtilsTrajectory {
    int32_t findNearestIndex(
        [in]  PLType("heapless::Vec<TrajectoryPoint, 10>")  points,
        [in]  PLType("nalgebra::Vector3<f64>")  query_position);
};

[generate(RustAWKPlugin, "")]
celltype tUtilsTrajectory {
    entry sUtilsTrajectory eUtils;
};