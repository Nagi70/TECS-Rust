import("struct_define.cdl");

signature sImuMsg {
};

signature sImuMsg {
};

signature sFrame {
};