import(<../spikert.cdl>);

cell tMotor Motor {
    port = C_EXP("PbioPortIdT::PbioPortIdA");
};

cell tSensor Sensor {
    port = C_EXP("PbioPortIdT::PbioPortIdC");
};

cell tMotorbody Motorbody {
    cMotor = Motor.eMotor;
};

cell tSensorbody Sensorbody {
    cSensor = Sensor.eSensor;
};

[generate( RustITRONPlugin, "lib, TASK")]
cell tTaskRs Task1{
    cTaskBody = Motorbody.eMotorbody;
    id = C_EXP("TECS_RUST_TASK1");
	task_ref = C_EXP("unsafe{TaskRef::from_raw_nonnull(NonZeroI32::new(TECS_RUST_TASK1).unwrap())}");
    attribute = C_EXP("TA_ACT");
    stackSize = 1024;
    priority = 7;
};

[generate( RustITRONPlugin, "lib, TASK")]
cell tTaskRs Task2{
    cTaskBody = Sensorbody.eSensorbody;
    id = C_EXP("TECS_RUST_TASK2");
	task_ref = C_EXP("unsafe{TaskRef::from_raw_nonnull(NonZeroI32::new(TECS_RUST_TASK2).unwrap())}");
    attribute = C_EXP("TA_ACT");
    stackSize = 1024;
    priority = 7;
};