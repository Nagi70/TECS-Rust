import("imu_driver.cdl");
import("awkernel_reactor.cdl");
import("diagnostic.cdl");

cell tReactor ImuReactor {
    cDagReactorbody = ImuDriver.eImuDriver;
    name = PL_EXP("imu_driver");
    schedType = PL_EXP("FIFO");
    publishTopicNames = PL_EXP("imu_raw");
    subscribeTopicNames = PL_EXP("imu");
    period = PL_EXP("Duration::from_sec(1)");
};

cell tImuDriver ImuDriver {
    cImuDriverbody = ImuDriverbody.eImuDriverbody;
};

cell tImuDriverbody ImuDriverbody {
    cDev      = ImuDev.eImuDevice;
    cRate     = RateMonitor.eRate;
    //period_ms = 5;
};

cell tTamagawaImuDevice ImuDev {
    can_id_gyro  = 0x319;
    can_id_accel = 0x31A;
    imu_frame_id = PL_EXP("imu");
};

cell tRateBoundStatus RateMonitor {
    reference_hz         = 200.0;
    ok_min_hz            = 100.0;
    ok_max_hz            = 10000.0;
    warn_min_hz          = 50.0;
    warn_max_hz          = 100000.0;
    num_frame_transition = 2;
};