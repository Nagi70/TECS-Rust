import("dummy_periodic_reactor.cdl");
import("publish_signature.cdl");
import("imu_driver.cdl");
import("imu_corrector.cdl");
import("vehicle_velocity_converter.cdl");
import("gyro_odometer.cdl");
import("ekf_localizer.cdl");

import("idx.cdl");

// IMU -> Ekf まで

cell tDummyPeriodicReactorInMrm DummyHardware {
    cImu = ImuDriver.eImu;
    cVelocityStatus = VehicleVelocityConverter.eVelocityStatus;
};

cell tImuDriver ImuDriver {
    cImuRaw = ImuCorrector.eImuRaw;
    cDev = TamagawaCan.eImuDevice;
};

cell tTamagawaImuDevice TamagawaCan {
    can_id_gyro  = 0x319;
    can_id_accel = 0x31A;
};

cell tImuCorrector ImuCorrector {
    cImuData = GyroOdometer.eImuData;
    cTf = ImuCorrectorTf.eTf;
};

cell tTf ImuCorrectorTf {
    transform = PL_EXP("nalgebra::Quaternion::new(1.0, 2.0, 1.0, 2.0)");
};

cell tVehicleVelocityConverter VehicleVelocityConverter {
    cTwistWithCovarianceV = GyroOdometer.eTwistWithCovarianceV;
};

cell tGyroOdometer GyroOdometer {
    cTwistWithCovarianceG = EkfLocalizer.eTwistWithCovarianceG;
    cTf = GyroOdometerTf.eTf;
};

cell tTf GyroOdometerTf {
    transform = PL_EXP("nalgebra::Quaternion::new(2.0, 1.0, 2.0, 1.0)");
};

cell tEkfLocalizer EkfLocalizer {
    cTwistWithCovarianceQueue = TwistWithCovarianceQueue.eSet;
};

cell tTwistWithCovarianceAgedObjectQueue TwistWithCovarianceQueue {
};

// Ekf から trajectory_follower まで

import("covariance.cdl");
import("time_delay_kalman_filter.cdl");
import("mahalanobis.cdl");
import("measurement.cdl");
import("state_transition.cdl");
import("utils_geometry.cdl");

import("stop_filter.cdl");
import("twist2accel.cdl");
import("trajectory_follower.cdl");
import("utils_trajectory.cdl");
import("utils_pose_deviation.cdl");
import("dummy_sink_reactor.cdl");

cell tEkfLocalizerTimer EkfLocalizerTimer {
    cKinematicState[0] = StopFilter.eKinematicState;
    cKinematicState[1] = Twist2Accel.eKinematicState;

    cEkfModule = EkfModule.eEkfModule;
    cQueue = TwistWithCovarianceQueue.eGet;
};

cell tEkfModule EkfModule {
    cKalman = TimeDelayKalmanFilter.eKalman;
    cState = StateTransition.eState;
    cMeasure = Measurement.eMeasure;
    cMaha = Mahalanobis.eMaha;
    cCov = Covariance.eCov;
    cUtils = UtilsGeometry.eUtils;
};

cell tTimeDelayKalmanFilter TimeDelayKalmanFilter {
};

cell tStateTransition StateTransition {
};

cell tMeasurement Measurement {
};

cell tMahalanobis Mahalanobis {
};

cell tCovariance Covariance {
};

cell tUtilsGeometry UtilsGeometry {
};

cell tStopFilter StopFilter {
    cKinematicStateSf = TrajectoryFollower.eKinematicStateSf;
};

cell tTwist2Accel Twist2Accel {
    cAccel = TrajectoryFollower.eAccel;
    
    cFilterAlx = FilterAlx.eFilter;
    cFilterAly = FilterAly.eFilter;
    cFilterAlz = FilterAlz.eFilter;
    cFilterAax = FilterAax.eFilter;
    cFilterAay = FilterAay.eFilter;
    cFilterAaz = FilterAaz.eFilter;
};

cell tLowpassFilter1D FilterAlx{
};

cell tLowpassFilter1D FilterAly{
};

cell tLowpassFilter1D FilterAlz{
};

cell tLowpassFilter1D FilterAax{
};

cell tLowpassFilter1D FilterAay{
};

cell tLowpassFilter1D FilterAaz{
};

cell tTrajectoryFollower TrajectoryFollower {
    cTraj = UtilsTrajectory.eUtils;
    cPose = UtilsPoseDeviation.eUtils;
    cControl = DummySinkReactor.eControl;
};

cell tUtilsTrajectory UtilsTrajectory {
};

cell tUtilsPoseDeviation UtilsPoseDeviation {
};

cell tDummySinkReactorInMrm DummySinkReactor {  
};