import("struct_define.cdl");
import("topic_signature.cdl");

signature sDummyImubody{
    void main([out] struct Frame* imu);
};

signature sDummyImuCorrectorbody{
    void main([in] struct ImuMsg imu_raw);
};

[generate( RustAWKPlugin, "")]
celltype tDummyImu{
    [async] call sDummyImubody cDummyImubody;
    entry sReactorbody eDummyImu;
};

[generate( RustAWKPlugin, "")]
celltype tDummyImuCorrector{
    [async] call sDummyImuCorrectorbody cDummyImuCorrectorbody;
    entry sReactorbody eDummyImuCorrector;
};

[generate( RustAWKPlugin, "")]
celltype tDummyImubody{
    [omit] call sImu cImu;
    entry sDummyImubody eDummyImubody;
};

[generate( RustAWKPlugin, "")]
celltype tDummyImuCorrectorbody{
    entry sImuRaw eImuRaw;
    entry sDummyImuCorrectorbody eDummyImuCorrectorbody;
};