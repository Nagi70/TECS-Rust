signature sArray {
    void main( [in] int32_t value );
};

signature sArrayTest {
    void main( [out] int32_t *value);
};

signature sInt {
    void send( [in] int32_t value);
};

[generate(RustAWKPlugin, "DAG_PERIODIC_REACTOR_BODY")]
celltype tArrayTest {
    call sArray cArray1;
    call sArray cArray2;

    entry sArrayTest eReactor;

    [omit] call sInt cInt;

    attr{
	    [omit] PLType("Cow") reactorName  = PL_EXP("ArrayTest");
	    [omit] PLType("SchedulerType") schedType = PL_EXP("SchedulerType::PrioritizedFIFO(7)");
	    [omit] PLType("Duration") period = PL_EXP("Duration::from_millis(50)");
        [omit] PLType("Cow") publishTopicNames = PL_EXP("Int");
    };
};

signature sDummy {
    void main( [in] int32_t value);
};

[generate(RustAWKPlugin, "DAG_SINK_REACTOR_BODY")]
celltype tDummy {
    entry sDummy eReactor;

    entry sInt eInt;

    attr{
	    [omit] PLType("Cow") reactorName  = PL_EXP("Dummy");
	    [omit] PLType("SchedulerType") schedType = PL_EXP("SchedulerType::PrioritizedFIFO(7)");
        [omit] PLType("Cow") subscribeTopicNames = PL_EXP("Int");
        [omit] PLType("Duration") relativeDeadline = PL_EXP("Duration::from_secs(1)");
    };
};

[generate(RustAWKPlugin, "")]
celltype tArray {

    entry sArray eArray;

  attr {
    [omit] int32_t  array_size = 2;

    [size_is(array_size)]
    int32_t  *attr_array;
  };
  var {
    [size_is(array_size)]
    int32_t  *var_array;
  };
};

cell tArrayTest ArrayTest {
    cArray1 = Array1.eArray;
    cArray2 = Array2.eArray;

    cInt = Dummy.eInt;
};

cell tDummy Dummy {
};

cell tArray Array1 {
    array_size = 1;
    attr_array = { 0 };
};

cell tArray Array2 {
    array_size = 2;
    attr_array = { 0, 0 };
};