import(<PaperSampleCelltype.cdl>);

[generate( RustITRONPlugin, "lib")]
cell tTaskRs Task1{
    cTaskBody = Manager.eManage1;
    id = C_EXP("TASK1");
	task_ref = C_EXP("unsafe{TaskRef::from_raw_nonnull(NonZeroI32::new(TASK1).unwrap())}");
    attribute = C_EXP("TA_ACT");
    stackSize = 1024;
    priority = 42;
};

[generate( RustITRONPlugin, "lib")]
cell tTaskRs Task2{
    cTaskBody = Taskbody1.eTaskbody;
    id = C_EXP("TASK2");
	task_ref = C_EXP("unsafe{TaskRef::from_raw_nonnull(NonZeroI32::new(TASK2).unwrap())}");
    attribute = C_EXP("TA_ACT");
    stackSize = 1024;
    priority = 42;
};

[generate( RustITRONPlugin, "lib")]
cell tTaskRs Task3{
    cTaskBody = Taskbody2.eTaskbody;
    id = C_EXP("TASK3");
	task_ref = C_EXP("unsafe{TaskRef::from_raw_nonnull(NonZeroI32::new(TASK3).unwrap())}");
    attribute = C_EXP("TA_ACT");
    stackSize = 1024;
    priority = 42;
};

cell tTaskbody1 Taskbody1 {
    cMotor = Motor2.eMotor;
    cManager = Manager.eManage2;
};

cell tManager Manager {
    cMotor = Motor1.eMotor;
};

cell tTaskbody2 Taskbody2 {
    cMotor = Motor2.eMotor;
    cSensor = Sensor.eSensor;
};

cell tMotor Motor1 {
    port = C_EXP("pbio_port_id_t::PBIO_PORT_ID_A");
};

cell tMotor Motor2 {
    port = C_EXP("pbio_port_id_t::PBIO_PORT_ID_B");
};

cell tSensor Sensor {
    port = C_EXP("pbio_port_id_t::PBIO_PORT_ID_C");
};
