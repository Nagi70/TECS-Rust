signature sHello {
    void hello(void);
};

signature sHello2 {
    void hello2(void);
};

signature sHello3 {
    void hello3(void);
};


signature sTaskbody {
    void main(void);
};

[active]
celltype tTask{
    call sTaskbody cTaskbody;
    attr {
        int32_t id;
    };
};

[generate(ItronrsGenPlugin,"lib")]
celltype tTaskbody {
    call sHello cPerson;
    entry sTaskbody eTaskbody;
};

[generate(ItronrsGenPlugin,"lib")]
celltype tAlice {
    call sHello2 cBob;
    call sHello2 cBob2;
    entry sHello eAlice1;
    entry sHello eAlice2;
    attr{
        int32_t id;
    };

    var{
        int32_t count = 0;
    };
};

[generate(ItronrsGenPlugin,"lib")]
celltype tBob {
    call sHello3 cCarol;
    entry sHello2 eBob1;
    entry sHello eBob2;
    attr{
        int32_t id;
    };

    var{
        int32_t count = 0;
    };
};

[generate(ItronrsGenPlugin,"lib")]
celltype tCarol {
    entry sHello3 eCarol;
    attr{
        int32_t id;
    };

    var{
        int32_t count = 0;
    };
};

[generate(ItronrsGenPlugin,"lib")]
cell tTask Task1 {
    cTaskbody = Taskbody1.eTaskbody;
    id = 0;
};

[generate(ItronrsGenPlugin,"lib")]
cell tTask Task2 {
    cTaskbody = Taskbody2.eTaskbody;
    id = 0;
};

[generate(ItronrsGenPlugin,"lib")]
cell tTask Task3 {
    cTaskbody = Taskbody3.eTaskbody;
    id = 0;
};

cell tTaskbody Taskbody1 {
    cPerson = Alice.eAlice1;
};

cell tTaskbody Taskbody2 {
    cPerson = Alice.eAlice2;
};

cell tTaskbody Taskbody3 {
    cPerson = Bob2.eBob2;
};

cell tAlice Alice {
    cBob = Bob.eBob1;
    cBob2 = Bob2.eBob1;
    id = 0;
};

cell tBob Bob {
    cCarol = Carol.eCarol;
    id = 1;
};

cell tBob Bob2 {
    cCarol = Carol2.eCarol;
    id = 2;
};

cell tCarol Carol {
    id = 1;
};

cell tCarol Carol2 {
    id = 2;
};