struct Header {
    PLType("awkernel_lib::time::Time") time_stamp;
    [string(256)] char* frame_id;
};

struct Frame {
    struct Header header;
    uint32_t id;
    bool_t is_rtr;
    bool_t is_extended;
    bool_t is_error;
    uint8_t dlc;
    uint8_t data[8];
};

struct ImuMsg {
    struct Header header;

    PLType("nalgebra::Quaternion<f64>")    orientation;                    /* geometry_msgs/Quaternion        */
    PLType("nalgebra::Matrix3<f64>")       orientation_covariance;

    PLType("nalgebra::Vector3<f64>")       angular_velocity;               /* geometry_msgs/Vector3           */
    PLType("nalgebra::Matrix3<f64>")       angular_velocity_covariance;

    PLType("nalgebra::Vector3<f64>")       linear_acceleration;            /* geometry_msgs/Vector3           */
    PLType("nalgebra::Matrix3<f64>")       linear_acceleration_covariance;
};

struct Twist {
    PLType("nalgebra::Vector3<f64>") linear;
    PLType("nalgebra::Vector3<f64>") angular;
};

struct TwistStamped {
    struct Header header;
    struct Twist twist;
};

struct TwistWithCovariance {
    struct Twist twist;           /* Twist 本体                           */
    PLType("nalgebra::Matrix6<f64>")       covariance;  /* 6x6 行列を 1 次元に展開               */
};

struct TwistWithCovarianceStamped {
    struct Header header;
    struct TwistWithCovariance      twist;      /* Twist + Covariance         */
};

struct VelocityReport {
    struct Header header;
    float32_t longitudinal_velocity;
    float32_t lateral_velocity;
    float32_t heading_rate;
};

struct Pose {
    PLType("nalgebra::Vector3<f64>")    point;
    PLType("nalgebra::Quaternion<f64>")    orientation;
};

struct PoseStamped {
    struct Header header;
    struct Pose      pose;      /* Twist + Covariance         */
};

struct PoseWithCovariance {
    struct Pose    pose;
    PLType("nalgebra::Matrix6<f64>")    covariance;
};

struct PoseWithCovarianceStamped {
    struct Header header;
    struct PoseWithCovariance      pose;      /* Twist + Covariance         */
};

struct Accel {
    PLType("nalgebra::Vector3<f64>") linear;
    PLType("nalgebra::Vector3<f64>") angular;
};

struct AccelWithCovariance {
    struct Accel    accel;
    PLType("nalgebra::Matrix6<f64>")    covariance;
};

struct AccelWithCovarianceStamped {
    struct Header header;
    struct AccelWithCovariance      accel;      /* Twist + Covariance         */
};

struct KinematicState {
    struct Header header;
    [string(256)] char* child_frame_id;
    struct PoseWithCovariance pose;
    struct TwistWithCovariance twist;
    struct AccelWithCovariance accel;
};

struct Transform {
    PLType("nalgebra::Vector3<f64>") translation;
    PLType("nalgebra::Quaternion<f64>") rotation;
};

/* Trajectory（autoware_planning_msgs/Trajectory の最小部分） */
struct TrajectoryPoint {
    struct Pose pose;
    double64_t longitudinal_velocity_mps;
};

/* TECS では可変長配列は PLType で表現。容量は固定（例: 5000点） */
struct Trajectory {
    struct Header header;
    PLType("heapless::Vec<TrajectoryPoint, 5000>") points;
};

struct Lateral {
    PLType("awkernel_lib::time::Time") stamp;
    double64_t steering_tire_angle;
};

struct Longitudinal {
    PLType("awkernel_lib::time::Time") stamp;
    double64_t velocity;
    double64_t acceleration;
};

struct Control {
    PLType("awkernel_lib::time::Time") stamp;
    struct Lateral lateral;
    struct Longitudinal longitudinal;
};