signature sHello {
    void hello(void);
};

signature sTaskbody {
    void main(void);
};

[active]
celltype tTask{
    call sTaskbody cTaskbody;
    attr {
        int32_t id;
    };
};

[generate(ItronrsGenPlugin,"lib")]
celltype tTaskbody {
    call sHello cPerson;
    entry sTaskbody eTaskbody;
};

[generate(ItronrsGenPlugin,"lib")]
celltype tAlice {
    call sHello cBob;
    entry sHello eAlice1;
    entry sHello eAlice2;
    entry sHello eAlice3;
    attr{
        int32_t id;
    };

    var{
        int32_t count = 0;
    };
};

[generate(ItronrsGenPlugin,"lib")]
celltype tBob {
    call sHello cAlice;
    entry sHello eBob;
    attr{
        int32_t id;
    };

    var{
        int32_t count = 0;
    };
};

[generate(ItronrsGenPlugin,"lib")]
cell tTask Task1 {
    cTaskbody = Taskbody1.eTaskbody;
    id = 0;
};

[generate(ItronrsGenPlugin,"lib")]
cell tTask Task2 {
    cTaskbody = Taskbody2.eTaskbody;
    id = 0;
};

cell tTaskbody Taskbody1 {
    cPerson = Alice.eAlice1;
};

cell tTaskbody Taskbody2 {
    cPerson = Alice.eAlice2;
};

cell tAlice Alice {
    cBob = Bob.eBob;
    id = 0;
};

cell tBob Bob {
    cAlice = Alice.eAlice3;
    id = 0;
};