import(<kernel_rs.cdl>);

typedef int_t   pbio_direction_t;
typedef int_t   pbio_port_id_t;
typedef int_t   pbio_error_t;
typedef int_t   Option_Ref_a_mut__pup_motor_t__;
typedef int_t   Option_Ref_a_mut__pup_ultrasonic_sensor_t__;
typedef int_t   bool;

signature sMotor {
    void set_motor_ref( void );
    void setup( [in] pbio_direction_t positive_direction, [in] bool reset_count );
    void set_speed( [in] int32_t speed );
    void stop( void );
};

signature sSensor {
    void set_device_ref( void );
    void get_distance( [out] int32_t* distance );
    void light_on( void );
    void light_set( [in] int32_t bv1, [in] int32_t bv2, [in] int32_t bv3, [in] int32_t bv4 );
    void light_off( void );
};

signature sPowerdown{
    void powerdown( [in] pbio_error_t error );
};

[generate (RustGenPlugin, "lib")]
celltype tMotor {
    call sPowerdown cPowerdown;
    [inline] entry sMotor eMotor;
    attr {
        pbio_port_id_t port = C_EXP("pbio_port_id_t::PBIO_PORT_ID_$port$");
    };
    var {
       Option_Ref_a_mut__pup_motor_t__ motor = C_EXP("None");
    };
};

[generate (RustGenPlugin, "lib")]
celltype tSensor {
    call sPowerdown cPowerdown;
    [inline] entry sSensor eSensor;
    attr{
        pbio_port_id_t port = C_EXP("pbio_port_id_t::PBIO_PORT_ID_$port$");
    };
    var {
        // RS_EXPもしくは，両方，もしくは別の表現，NONTECS_EXPみたいな
        Option_Ref_a_mut__pup_ultrasonic_sensor_t__ ult = C_EXP("None");
    };
};

[generate (RustGenPlugin, "lib")]
celltype tTaskbody {
    [inline] entry sTaskBody eTaskbody;
    call sSensor cSensor;
    call sMotor cMotor;
};

[generate (RustGenPlugin, "lib")]
celltype tPowerdown {
    [inline] entry sPowerdown ePowerdown1;
    [inline] entry sPowerdown ePowerdown2;
};

cell tMotor Motor {
    cPowerdown = Powerdown.ePowerdown1;
    port = C_EXP("pbio_port_id_t::PBIO_PORT_ID_A");
};

cell tSensor Sensor {
    cPowerdown = Powerdown.ePowerdown2;
    port = C_EXP("pbio_port_id_t::PBIO_PORT_ID_B");
};

cell tTaskbody Taskbody {
    cMotor = Motor.eMotor;
    cSensor = Sensor.eSensor;
};

cell tPowerdown Powerdown{
};

[generate( RustITRONPlugin, "lib")]
cell tTask_rs Task{
    cTaskBody = Taskbody.eTaskbody;
    id = C_EXP("TASK1");
	task_ref = C_EXP("unsafe{TaskRef::from_raw_nonnull(NonZeroI32::new(TASK1).unwrap())}");
    attribute = C_EXP("TA_ACT");
    stackSize = 1024;
    priority = 42;
};