struct ImuData {
    RType("Time")     time_stamp;                /* [us] */
    float32_t    angular_velocity_x;        /* [rad/s] */
    float32_t    angular_velocity_y;        /* [rad/s] */
    float32_t    angular_velocity_z;        /* [rad/s] */
    float32_t    linear_acceleration_x;     /* [m/s^2] */
    float32_t    linear_acceleration_y;     /* [m/s^2] */
    float32_t    linear_acceleration_z;     /* [m/s^2] */
};

struct Header {
    RType("Time") time_stamp;
    [string(256)] char* frame_id;
};

struct Quaternion {
    double64_t x;
    double64_t y;
    double64_t z;
    double64_t w;
};

struct Vector3 {
    double64_t x;
    double64_t y;
    double64_t z;
};

struct ImuMsg {
    struct Header header;

    struct Quaternion    orientation;                    /* geometry_msgs/Quaternion        */
    double64_t        orientation_covariance[9];

    struct Vector3       angular_velocity;               /* geometry_msgs/Vector3           */
    double64_t        angular_velocity_covariance[9];

    struct Vector3       linear_acceleration;            /* geometry_msgs/Vector3           */
    double64_t        linear_acceleration_covariance[9];
};

struct Transform {
    struct Vector3    translation;                /* TF translation */
    struct Quaternion rotation;                   /* TF rotation    */
};

struct Twist {
    struct Vector3 linear;
    struct Vector3 angular;
};

struct TwistStamped {
    uint64_t time_stamp;          /* Header.stamp の代替 [ns]            */
    char_t  *frame_id;            /* Header.frame_id の代替               */
    struct Twist twist;           /* geometry_msgs/Twist                  */
};

struct TwistWithCovariance {
    struct Twist twist;           /* Twist 本体                           */
    double64_t       covariance[36];  /* 6x6 行列を 1 次元に展開               */
};

struct TwistWithCovarianceStamped {
    uint64_t                        time_stamp;  /* Header.stamp [ns]          */
    char_t                        *frame_id;    /* Header.frame_id            */
    struct TwistWithCovariance      twist;      /* Twist + Covariance         */
};

struct Frame {
    struct Header header;
    uint32_t id;
    bool_t is_rtr;
    bool_t is_extended;
    bool_t is_error;
    uint8_t dlc;
    uint8_t data[8];
};