signature sStateTransition {
    double64_t normalizeYaw( [in] double64_t yaw );
    PLType("nalgebra::Vector6<f64>") predictNextState( 
        [in] PLType("nalgebra::Vector6<f64>") x_curr,
        [in] double64_t dt
    );
    PLType("nalgebra::Matrix6<f64>") createStateTransitionMatrix( 
        [in] PLType("nalgebra::Vector6<f64>") x_curr,
        [in] double64_t dt
    );
    PLType("nalgebra::Matrix6<f64>") processNoiseCovariance( 
        [in] double64_t proc_cov_yaw_d,
        [in] double64_t proc_cov_vx_d,
        [in] double64_t proc_cov_wz_d
    );
};

[generate( RustAWKPlugin, "")]
celltype tStateTransition {
    entry sStateTransition eState;  
};